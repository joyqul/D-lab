module ELEVATOR(FLOOR, OPEN, CLK, RESET, PEOPLE, GOTO);

    input            CLK, RESET, PEOPLE; 
    input      [2:0] GOTO;
    output reg       OPEN;   
    output reg [2:0] FLOOR;






endmodule
